library ieee;
use ieee.std_logic_1164.all;


entity datapath is
    port(

    );
end datapath;

architecture logic of datapath is
begin
    
end logic;